--helloo
-- hello again
-- helloooooo