--helloo
